// Code your testbench here
// or browse Examples
//`include "memory_tb.sv"
//`include "regfile_tb.sv"
//`include "ALU_tb.sv"

//`include "risc_instructions_handler.sv"
//`include "test_code_tb.sv"

//`include "risc_instructions_handler_tb.sv"

`include "risc_v_tb.sv"



